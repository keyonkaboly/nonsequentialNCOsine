module test1;
  
  reg[15:0] regs[0:255];
  reg[15:0] opt;  
integer i;

initial begin
regs[0] = 0;
regs[1] = 804;
regs[2] = 1608;
regs[3] = 2410;
regs[4] = 3212;
regs[5] = 4011;
regs[6] = 4808;
regs[7] = 5602;
regs[8] = 6393;
regs[9] = 7179;
regs[10] = 7962;
regs[11] = 8739;
regs[12] = 9512;
regs[13] = 10278;
regs[14] = 11039;
regs[15] = 11793;
regs[16] = 12539;
regs[17] = 13279;
regs[18] = 14010;
regs[19] = 14732;
regs[20] = 15446;
regs[21] = 16151;
regs[22] = 16846;
regs[23] = 17530;
regs[24] = 18204;
regs[25] = 18868;
regs[26] = 19519;
regs[27] = 20159;
regs[28] = 20787;
regs[29] = 21403;
regs[30] = 22005;
regs[31] = 22594;
regs[32] = 23170;
regs[33] = 23731;
regs[34] = 24279;
regs[35] = 24811;
regs[36] = 25329;
regs[37] = 25832;
regs[38] = 26319;
regs[39] = 26790;
regs[40] = 27245;
regs[41] = 27683;
regs[42] = 28105;
regs[43] = 28510;
regs[44] = 28898;
regs[45] = 29268;
regs[46] = 29621;
regs[47] = 29956;
regs[48] = 30273;
regs[49] = 30571;
regs[50] = 30852;
regs[51] = 31113;
regs[52] = 31356;
regs[53] = 31580;
regs[54] = 31785;
regs[55] = 31971;
regs[56] = 32137;
regs[57] = 32285;
regs[58] = 32412;
regs[59] = 32521;
regs[60] = 32609;
regs[61] = 32678;
regs[62] = 32728;
regs[63] = 32757;
regs[64] = 32767;
regs[65] = 32757;
regs[66] = 32728;
regs[67] = 32678;
regs[68] = 32609;
regs[69] = 32521;
regs[70] = 32412;
regs[71] = 32285;
regs[72] = 32137;
regs[73] = 31971;
regs[74] = 31785;
regs[75] = 31580;
regs[76] = 31356;
regs[77] = 31113;
regs[78] = 30852;
regs[79] = 30571;
regs[80] = 30273;
regs[81] = 29956;
regs[82] = 29621;
regs[83] = 29268;
regs[84] = 28898;
regs[85] = 28510;
regs[86] = 28105;
regs[87] = 27683;
regs[88] = 27245;
regs[89] = 26790;
regs[90] = 26319;
regs[91] = 25832;
regs[92] = 25329;
regs[93] = 24811;
regs[94] = 24279;
regs[95] = 23731;
regs[96] = 23170;
regs[97] = 22594;
regs[98] = 22005;
regs[99] = 21403;
regs[100] = 20787;
regs[101] = 20159;
regs[102] = 19519;
regs[103] = 18868;
regs[104] = 18204;
regs[105] = 17530;
regs[106] = 16846;
regs[107] = 16151;
regs[108] = 15446;
regs[109] = 14732;
regs[110] = 14010;
regs[111] = 13279;
regs[112] = 12539;
regs[113] = 11793;
regs[114] = 11039;
regs[115] = 10278;
regs[116] = 9512;
regs[117] = 8739;
regs[118] = 7962;
regs[119] = 7179;
regs[120] = 6393;
regs[121] = 5602;
regs[122] = 4808;
regs[123] = 4011;
regs[124] = 3212;
regs[125] = 2410;
regs[126] = 1608;
regs[127] = 804;
regs[128] = 0;
regs[129] = -804;
regs[130] = -1608;
regs[131] = -2410;
regs[132] = -3212;
regs[133] = -4011;
regs[134] = -4808;
regs[135] = -5602;
regs[136] = -6393;
regs[137] = -7179;
regs[138] = -7962;
regs[139] = -8739;
regs[140] = -9512;
regs[141] = -10278;
regs[142] = -11039;
regs[143] = -11793;
regs[144] = -12539;
regs[145] = -13279;
regs[146] = -14010;
regs[147] = -14732;
regs[148] = -15446;
regs[149] = -16151;
regs[150] = -16846;
regs[151] = -17530;
regs[152] = -18204;
regs[153] = -18868;
regs[154] = -19519;
regs[155] = -20159;
regs[156] = -20787;
regs[157] = -21403;
regs[158] = -22005;
regs[159] = -22594;
regs[160] = -23170;
regs[161] = -23731;
regs[162] = -24279;
regs[163] = -24811;
regs[164] = -25329;
regs[165] = -25832;
regs[166] = -26319;
regs[167] = -26790;
regs[168] = -27245;
regs[169] = -27683;
regs[170] = -28105;
regs[171] = -28510;
regs[172] = -28898;
regs[173] = -29268;
regs[174] = -29621;
regs[175] = -29956;
regs[176] = -30273;
regs[177] = -30571;
regs[178] = -30852;
regs[179] = -31113;
regs[180] = -31356;
regs[181] = -31580;
regs[182] = -31785;
regs[183] = -31971;
regs[184] = -32137;
regs[185] = -32285;
regs[186] = -32412;
regs[187] = -32521;
regs[188] = -32609;
regs[189] = -32678;
regs[190] = -32728;
regs[191] = -32757;
regs[192] = -32767;
regs[193] = -32757;
regs[194] = -32728;
regs[195] = -32678;
regs[196] = -32609;
regs[197] = -32521;
regs[198] = -32412;
regs[199] = -32285;
regs[200] = -32137;
regs[201] = -31971;
regs[202] = -31785;
regs[203] = -31580;
regs[204] = -31356;
regs[205] = -31113;
regs[206] = -30852;
regs[207] = -30571;
regs[208] = -30273;
regs[209] = -29956;
regs[210] = -29621;
regs[211] = -29268;
regs[212] = -28898;
regs[213] = -28510;
regs[214] = -28105;
regs[215] = -27683;
regs[216] = -27245;
regs[217] = -26790;
regs[218] = -26319;
regs[219] = -25832;
regs[220] = -25329;
regs[221] = -24811;
regs[222] = -24279;
regs[223] = -23731;
regs[224] = -23170;
regs[225] = -22594;
regs[226] = -22005;
regs[227] = -21403;
regs[228] = -20787;
regs[229] = -20159;
regs[230] = -19519;
regs[231] = -18868;
regs[232] = -18204;
regs[233] = -17530;
regs[234] = -16846;
regs[235] = -16151;
regs[236] = -15446;
regs[237] = -14732;
regs[238] = -14010;
regs[239] = -13279;
regs[240] = -12539;
regs[241] = -11793;
regs[242] = -11039;
regs[243] = -10278;
regs[244] = -9512;
regs[245] = -8739;
regs[246] = -7962;
regs[247] = -7179;
regs[248] = -6393;
regs[249] = -5602;
regs[250] = -4808;
regs[251] = -4011;
regs[252] = -3212;
regs[253] = -2410;
regs[254] = -1608;
regs[255] = -804;

    for (i = 0; i < 256; i = i + 1) begin
      opt = regs[i];
      #20; 
    end
 
end

  initial begin
    $monitor("%0t .. %d", $time, opt);
  end
endmodule
